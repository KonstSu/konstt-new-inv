magic
tech sky130A
magscale 1 2
timestamp 1761058134
<< error_s >>
rect 2130 -100 2290 -96
rect 2600 -190 2676 -62
rect 2730 -100 4730 -96
rect 2718 -130 2720 -118
rect 4740 -130 4742 -118
rect 2730 -142 2742 -140
rect 4718 -142 4730 -140
rect 2182 -200 2240 -194
rect 2600 -196 4680 -190
rect 2182 -234 2194 -200
rect 2182 -240 2240 -234
rect 2336 -510 2422 -256
rect 2600 -402 2676 -196
rect 4540 -348 4541 -288
rect 4568 -376 4569 -281
rect 2590 -570 2676 -402
rect 2600 -700 2676 -570
rect 2182 -1528 2240 -1522
rect 2182 -1562 2194 -1528
rect 2182 -1568 2240 -1562
<< nwell >>
rect 4539 -349 4543 -284
rect 2590 -570 4590 -510
<< pwell >>
rect 4550 -1260 4680 -1210
rect 2700 -1550 4410 -1520
<< viali >>
rect 2130 -130 2290 -100
rect 2730 -130 4730 -100
rect 2130 -1670 2300 -1630
rect 2930 -1680 4560 -1640
<< metal1 >>
rect 1840 100 5000 500
rect 1840 -280 1980 100
rect 2100 -100 2320 100
rect 2100 -130 2130 -100
rect 2290 -130 2320 -100
rect 2100 -160 2320 -130
rect 2720 -100 4740 100
rect 2720 -130 2730 -100
rect 4730 -130 4740 -100
rect 2720 -140 4740 -130
rect 2510 -240 4680 -190
rect 2510 -280 2590 -240
rect 1840 -480 2180 -280
rect 2230 -480 2590 -280
rect 2727 -348 2737 -288
rect 2794 -348 2804 -288
rect 2920 -348 2930 -288
rect 2987 -348 2997 -288
rect 3113 -348 3123 -288
rect 3180 -348 3190 -288
rect 3306 -348 3316 -288
rect 3373 -348 3383 -288
rect 3499 -348 3509 -288
rect 3566 -348 3576 -288
rect 3692 -348 3702 -288
rect 3759 -348 3769 -288
rect 3885 -348 3895 -288
rect 3952 -348 3962 -288
rect 4078 -348 4088 -288
rect 4145 -348 4155 -288
rect 4271 -348 4281 -288
rect 4338 -348 4348 -288
rect 4464 -348 4474 -288
rect 4531 -348 4541 -288
rect 2460 -510 2590 -480
rect 1880 -570 2250 -520
rect 2460 -570 4590 -510
rect 1880 -800 1940 -570
rect 1500 -1000 1940 -800
rect 1880 -1220 1940 -1000
rect 2460 -1210 2590 -570
rect 5200 -1000 5400 -800
rect 1880 -1260 2260 -1220
rect 2460 -1260 4680 -1210
rect 2460 -1300 2590 -1260
rect 1880 -1480 2180 -1320
rect 2230 -1480 2590 -1300
rect 1880 -1900 2000 -1480
rect 2510 -1520 2590 -1480
rect 2510 -1560 4590 -1520
rect 2110 -1630 2320 -1610
rect 2110 -1670 2130 -1630
rect 2300 -1670 2320 -1630
rect 2110 -1680 2320 -1670
rect 2120 -1900 2320 -1680
rect 2720 -1640 4730 -1630
rect 2720 -1680 2930 -1640
rect 4560 -1680 4730 -1640
rect 2720 -1900 4730 -1680
rect 1880 -2300 5000 -1900
<< via1 >>
rect 2737 -348 2794 -288
rect 2930 -348 2987 -288
rect 3123 -348 3180 -288
rect 3316 -348 3373 -288
rect 3509 -348 3566 -288
rect 3702 -348 3759 -288
rect 3895 -348 3952 -288
rect 4088 -348 4145 -288
rect 4281 -348 4338 -288
rect 4474 -348 4531 -288
<< metal2 >>
rect 2737 -280 2794 -278
rect 2930 -280 2987 -278
rect 3123 -280 3180 -278
rect 3316 -280 3373 -278
rect 3509 -280 3566 -278
rect 3702 -280 3759 -278
rect 3895 -280 3952 -278
rect 4088 -280 4145 -278
rect 4281 -280 4338 -278
rect 4474 -280 4531 -278
rect 2720 -288 6477 -280
rect 2720 -348 2737 -288
rect 2794 -348 2930 -288
rect 2987 -348 3123 -288
rect 3180 -348 3316 -288
rect 3373 -348 3509 -288
rect 3566 -348 3702 -288
rect 3759 -348 3895 -288
rect 3952 -348 4088 -288
rect 4145 -348 4281 -288
rect 4338 -348 4474 -288
rect 4531 -348 6477 -288
rect 2720 -350 6477 -348
rect 2737 -358 2794 -350
rect 2930 -358 2987 -350
rect 3123 -358 3180 -350
rect 3316 -358 3373 -350
rect 3509 -358 3566 -350
rect 3702 -358 3759 -350
rect 3895 -358 3952 -350
rect 4088 -358 4145 -350
rect 4281 -358 4338 -350
rect 4474 -358 4531 -350
rect 2720 -480 4870 -420
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1 ~/asic/konstt-new-inv/mag
timestamp 1761054031
transform 1 0 2211 0 -1 -381
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM2 ~/asic/konstt-new-inv/mag
timestamp 1761054031
transform 1 0 2211 0 1 -1390
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_8DVCWJ  XM3 ~/asic/konstt-new-inv/mag
timestamp 1761054031
transform 1 0 3727 0 1 -381
box -1127 -319 1127 319
use sky130_fd_pr__nfet_01v8_YTLFGX  XM4 ~/asic/konstt-new-inv/mag
timestamp 1761054031
transform 1 0 3727 0 1 -1390
box -1127 -310 1127 310
<< labels >>
flabel metal1 1500 -1000 1700 -800 0 FreeSans 256 0 0 0 in0
port 3 nsew
flabel metal1 5200 -1000 5400 -800 0 FreeSans 256 0 0 0 out0
port 2 nsew
flabel metal1 2100 200 2300 400 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 2100 -2200 2300 -2000 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
