magic
tech sky130A
magscale 1 2
timestamp 1758902349
<< error_s >>
rect 2130 -100 2300 -96
rect 2182 -200 2240 -194
rect 3082 -200 3140 -194
rect 3274 -200 3332 -194
rect 3466 -200 3524 -194
rect 3658 -200 3716 -194
rect 3850 -200 3908 -194
rect 4042 -200 4100 -194
rect 4234 -200 4292 -194
rect 4426 -200 4484 -194
rect 4618 -200 4676 -194
rect 4810 -200 4868 -194
rect 2182 -234 2194 -200
rect 3082 -234 3094 -200
rect 3274 -234 3286 -200
rect 3466 -234 3478 -200
rect 3658 -234 3670 -200
rect 3850 -234 3862 -200
rect 4042 -234 4054 -200
rect 4234 -234 4246 -200
rect 4426 -234 4438 -200
rect 4618 -234 4630 -200
rect 4810 -234 4822 -200
rect 2182 -240 2240 -234
rect 3082 -240 3140 -234
rect 3274 -240 3332 -234
rect 3466 -240 3524 -234
rect 3658 -240 3716 -234
rect 3850 -240 3908 -234
rect 4042 -240 4100 -234
rect 4234 -240 4292 -234
rect 4426 -240 4484 -234
rect 4618 -240 4676 -234
rect 4810 -240 4868 -234
rect 2182 -528 2240 -522
rect 2986 -528 3044 -522
rect 3178 -528 3236 -522
rect 3370 -528 3428 -522
rect 3562 -528 3620 -522
rect 3754 -528 3812 -522
rect 3946 -528 4004 -522
rect 4138 -528 4196 -522
rect 4330 -528 4388 -522
rect 4522 -528 4580 -522
rect 4714 -528 4772 -522
rect 2182 -562 2194 -528
rect 2986 -562 2998 -528
rect 3178 -562 3190 -528
rect 3370 -562 3382 -528
rect 3562 -562 3574 -528
rect 3754 -562 3766 -528
rect 3946 -562 3958 -528
rect 4138 -562 4150 -528
rect 4330 -562 4342 -528
rect 4522 -562 4534 -528
rect 4714 -562 4726 -528
rect 2182 -568 2240 -562
rect 2986 -568 3044 -562
rect 3178 -568 3236 -562
rect 3370 -568 3428 -562
rect 3562 -568 3620 -562
rect 3754 -568 3812 -562
rect 3946 -568 4004 -562
rect 4138 -568 4196 -562
rect 4330 -568 4388 -562
rect 4522 -568 4580 -562
rect 4714 -568 4772 -562
rect 2182 -1218 2240 -1212
rect 3082 -1218 3140 -1212
rect 3274 -1218 3332 -1212
rect 3466 -1218 3524 -1212
rect 3658 -1218 3716 -1212
rect 3850 -1218 3908 -1212
rect 4042 -1218 4100 -1212
rect 4234 -1218 4292 -1212
rect 4426 -1218 4484 -1212
rect 4618 -1218 4676 -1212
rect 4810 -1218 4868 -1212
rect 2182 -1252 2194 -1218
rect 3082 -1252 3094 -1218
rect 3274 -1252 3286 -1218
rect 3466 -1252 3478 -1218
rect 3658 -1252 3670 -1218
rect 3850 -1252 3862 -1218
rect 4042 -1252 4054 -1218
rect 4234 -1252 4246 -1218
rect 4426 -1252 4438 -1218
rect 4618 -1252 4630 -1218
rect 4810 -1252 4822 -1218
rect 2182 -1258 2240 -1252
rect 3082 -1258 3140 -1252
rect 3274 -1258 3332 -1252
rect 3466 -1258 3524 -1252
rect 3658 -1258 3716 -1252
rect 3850 -1258 3908 -1252
rect 4042 -1258 4100 -1252
rect 4234 -1258 4292 -1252
rect 4426 -1258 4484 -1252
rect 4618 -1258 4676 -1252
rect 4810 -1258 4868 -1252
rect 2182 -1528 2240 -1522
rect 2986 -1528 3044 -1522
rect 3178 -1528 3236 -1522
rect 3370 -1528 3428 -1522
rect 3562 -1528 3620 -1522
rect 3754 -1528 3812 -1522
rect 3946 -1528 4004 -1522
rect 4138 -1528 4196 -1522
rect 4330 -1528 4388 -1522
rect 4522 -1528 4580 -1522
rect 4714 -1528 4772 -1522
rect 2182 -1562 2194 -1528
rect 2986 -1562 2998 -1528
rect 3178 -1562 3190 -1528
rect 3370 -1562 3382 -1528
rect 3562 -1562 3574 -1528
rect 3754 -1562 3766 -1528
rect 3946 -1562 3958 -1528
rect 4138 -1562 4150 -1528
rect 4330 -1562 4342 -1528
rect 4522 -1562 4534 -1528
rect 4714 -1562 4726 -1528
rect 2182 -1568 2240 -1562
rect 2986 -1568 3044 -1562
rect 3178 -1568 3236 -1562
rect 3370 -1568 3428 -1562
rect 3562 -1568 3620 -1562
rect 3754 -1568 3812 -1562
rect 3946 -1568 4004 -1562
rect 4138 -1568 4196 -1562
rect 4330 -1568 4388 -1562
rect 4522 -1568 4580 -1562
rect 4714 -1568 4772 -1562
<< viali >>
rect 2130 -130 2300 -100
rect 2130 -1670 2300 -1630
<< metal1 >>
rect 2000 100 5000 500
rect 2100 -100 2320 100
rect 2100 -130 2130 -100
rect 2300 -130 2320 -100
rect 2100 -160 2320 -130
rect 1500 -1000 1700 -800
rect 5200 -1000 5400 -800
rect 2110 -1630 2320 -1610
rect 2110 -1670 2130 -1630
rect 2300 -1670 2320 -1630
rect 2110 -1680 2320 -1670
rect 2120 -1900 2320 -1680
rect 2000 -2300 5000 -1900
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1758902349
transform 1 0 2211 0 1 -381
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1758902349
transform 1 0 2211 0 1 -1390
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_8DVCWJ  XM3
timestamp 1758902349
transform 1 0 3927 0 1 -381
box -1127 -319 1127 319
use sky130_fd_pr__nfet_01v8_YTLFGX  XM4
timestamp 1758902349
transform 1 0 3927 0 1 -1390
box -1127 -310 1127 310
<< labels >>
flabel metal1 1500 -1000 1700 -800 0 FreeSans 256 0 0 0 in0
port 3 nsew
flabel metal1 5200 -1000 5400 -800 0 FreeSans 256 0 0 0 out0
port 2 nsew
flabel metal1 2100 200 2300 400 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 2100 -2200 2300 -2000 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
