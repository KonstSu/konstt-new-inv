magic
tech sky130A
magscale 1 2
timestamp 1761646426
<< nwell >>
rect 4390 70 4750 420
rect 2710 -250 4750 70
<< viali >>
rect 3180 -30 4350 30
rect 2010 -100 2140 -60
rect 2000 -1660 2130 -1620
rect 3180 -1700 4430 -1640
<< metal1 >>
rect 1760 380 4850 500
rect 1760 150 4430 380
rect 4700 150 4850 380
rect 1760 110 4850 150
rect 1760 -170 1840 110
rect 1980 -60 2160 110
rect 2700 70 4750 110
rect 2700 30 4730 70
rect 2700 -30 3180 30
rect 4350 -30 4730 30
rect 2700 -40 4730 -30
rect 1980 -100 2010 -60
rect 2140 -100 2160 -60
rect 1980 -110 2160 -100
rect 2340 -150 4670 -90
rect 2340 -170 2510 -150
rect 1760 -390 2050 -170
rect 2100 -380 2510 -170
rect 2710 -240 2720 -180
rect 2790 -240 2800 -180
rect 2910 -240 2920 -182
rect 2981 -240 2991 -182
rect 3099 -240 3109 -182
rect 3170 -240 3180 -182
rect 3293 -239 3303 -181
rect 3364 -239 3374 -181
rect 3483 -240 3493 -182
rect 3554 -240 3564 -182
rect 3676 -240 3686 -182
rect 3747 -240 3757 -182
rect 3867 -240 3877 -182
rect 3938 -240 3948 -182
rect 4062 -240 4072 -182
rect 4133 -240 4143 -182
rect 4252 -240 4262 -182
rect 4323 -240 4333 -182
rect 4444 -240 4454 -182
rect 4515 -240 4525 -182
rect 4637 -238 4647 -180
rect 4708 -238 4718 -180
rect 2812 -371 2822 -313
rect 2883 -371 2893 -313
rect 3005 -370 3015 -312
rect 3076 -370 3086 -312
rect 3196 -370 3206 -312
rect 3267 -370 3277 -312
rect 3387 -372 3397 -314
rect 3458 -372 3468 -314
rect 3581 -370 3591 -312
rect 3652 -370 3662 -312
rect 3775 -372 3785 -314
rect 3846 -372 3856 -314
rect 3964 -372 3974 -314
rect 4035 -372 4045 -314
rect 4157 -372 4167 -314
rect 4228 -372 4238 -314
rect 4348 -370 4358 -312
rect 4419 -370 4429 -312
rect 4540 -372 4550 -314
rect 4611 -372 4621 -314
rect 2340 -420 2510 -380
rect 1650 -510 2110 -420
rect 2340 -490 4580 -420
rect 1650 -800 1760 -510
rect 1420 -1000 1760 -800
rect 1650 -1230 1760 -1000
rect 2340 -1200 2510 -490
rect 4410 -810 5400 -800
rect 4410 -990 4420 -810
rect 4720 -990 5400 -810
rect 4410 -1000 5400 -990
rect 1650 -1310 2120 -1230
rect 2340 -1260 4650 -1200
rect 2340 -1340 2510 -1260
rect 1650 -1540 2040 -1340
rect 2100 -1520 2510 -1340
rect 2700 -1349 2710 -1289
rect 2780 -1349 2790 -1289
rect 2900 -1349 2910 -1291
rect 2971 -1349 2981 -1291
rect 3089 -1349 3099 -1291
rect 3160 -1349 3170 -1291
rect 3283 -1348 3293 -1290
rect 3354 -1348 3364 -1290
rect 3473 -1349 3483 -1291
rect 3544 -1349 3554 -1291
rect 3666 -1349 3676 -1291
rect 3737 -1349 3747 -1291
rect 3857 -1349 3867 -1291
rect 3928 -1349 3938 -1291
rect 4052 -1349 4062 -1291
rect 4123 -1349 4133 -1291
rect 4242 -1349 4252 -1291
rect 4313 -1349 4323 -1291
rect 4434 -1349 4444 -1291
rect 4505 -1349 4515 -1291
rect 4627 -1347 4637 -1289
rect 4698 -1347 4708 -1289
rect 2800 -1479 2810 -1421
rect 2871 -1479 2881 -1421
rect 2993 -1478 3003 -1420
rect 3064 -1478 3074 -1420
rect 3184 -1478 3194 -1420
rect 3255 -1478 3265 -1420
rect 3375 -1480 3385 -1422
rect 3446 -1480 3456 -1422
rect 3569 -1478 3579 -1420
rect 3640 -1478 3650 -1420
rect 3763 -1480 3773 -1422
rect 3834 -1480 3844 -1422
rect 3952 -1480 3962 -1422
rect 4023 -1480 4033 -1422
rect 4145 -1480 4155 -1422
rect 4216 -1480 4226 -1422
rect 4336 -1478 4346 -1420
rect 4407 -1478 4417 -1420
rect 4528 -1480 4538 -1422
rect 4599 -1480 4609 -1422
rect 2100 -1540 4560 -1520
rect 1650 -1940 1830 -1540
rect 2360 -1570 4560 -1540
rect 1980 -1620 2160 -1600
rect 1980 -1660 2000 -1620
rect 2130 -1660 2160 -1620
rect 1980 -1940 2160 -1660
rect 2690 -1640 4710 -1630
rect 2690 -1700 3180 -1640
rect 4430 -1700 4710 -1640
rect 2690 -1940 4710 -1700
rect 1650 -1950 4800 -1940
rect 1650 -2240 4360 -1950
rect 4680 -2240 4800 -1950
rect 1650 -2300 4800 -2240
<< via1 >>
rect 4430 150 4700 380
rect 2720 -240 2790 -180
rect 2920 -240 2981 -182
rect 3109 -240 3170 -182
rect 3303 -239 3364 -181
rect 3493 -240 3554 -182
rect 3686 -240 3747 -182
rect 3877 -240 3938 -182
rect 4072 -240 4133 -182
rect 4262 -240 4323 -182
rect 4454 -240 4515 -182
rect 4647 -238 4708 -180
rect 2822 -371 2883 -313
rect 3015 -370 3076 -312
rect 3206 -370 3267 -312
rect 3397 -372 3458 -314
rect 3591 -370 3652 -312
rect 3785 -372 3846 -314
rect 3974 -372 4035 -314
rect 4167 -372 4228 -314
rect 4358 -370 4419 -312
rect 4550 -372 4611 -314
rect 4420 -990 4720 -810
rect 2710 -1349 2780 -1289
rect 2910 -1349 2971 -1291
rect 3099 -1349 3160 -1291
rect 3293 -1348 3354 -1290
rect 3483 -1349 3544 -1291
rect 3676 -1349 3737 -1291
rect 3867 -1349 3928 -1291
rect 4062 -1349 4123 -1291
rect 4252 -1349 4313 -1291
rect 4444 -1349 4505 -1291
rect 4637 -1347 4698 -1289
rect 2810 -1479 2871 -1421
rect 3003 -1478 3064 -1420
rect 3194 -1478 3255 -1420
rect 3385 -1480 3446 -1422
rect 3579 -1478 3640 -1420
rect 3773 -1480 3834 -1422
rect 3962 -1480 4023 -1422
rect 4155 -1480 4216 -1422
rect 4346 -1478 4407 -1420
rect 4538 -1480 4599 -1422
rect 4360 -2240 4680 -1950
<< metal2 >>
rect 4390 380 4750 420
rect 4390 150 4430 380
rect 4700 150 4750 380
rect 4390 70 4750 150
rect 2710 -180 4750 70
rect 2710 -240 2720 -180
rect 2790 -181 4647 -180
rect 2790 -182 3303 -181
rect 2790 -240 2920 -182
rect 2981 -240 3109 -182
rect 3170 -239 3303 -182
rect 3364 -182 4647 -181
rect 3364 -239 3493 -182
rect 3170 -240 3493 -239
rect 3554 -240 3686 -182
rect 3747 -240 3877 -182
rect 3938 -240 4072 -182
rect 4133 -240 4262 -182
rect 4323 -240 4454 -182
rect 4515 -238 4647 -182
rect 4708 -238 4750 -180
rect 4515 -240 4750 -238
rect 2710 -250 4750 -240
rect 2822 -313 2883 -303
rect 2710 -371 2822 -320
rect 3015 -312 3076 -302
rect 2883 -370 3015 -320
rect 3206 -312 3267 -302
rect 3076 -370 3206 -320
rect 3397 -314 3458 -304
rect 3267 -370 3397 -320
rect 2883 -371 3397 -370
rect 2710 -372 3397 -371
rect 3591 -312 3652 -302
rect 3458 -370 3591 -320
rect 3785 -314 3846 -304
rect 3652 -370 3785 -320
rect 3458 -372 3785 -370
rect 3974 -314 4035 -304
rect 3846 -372 3974 -320
rect 4167 -314 4228 -304
rect 4035 -372 4167 -320
rect 4358 -312 4419 -302
rect 4228 -370 4358 -320
rect 4550 -314 4611 -304
rect 4419 -370 4550 -320
rect 4228 -372 4550 -370
rect 4611 -372 4740 -320
rect 2710 -620 4740 -372
rect 4390 -810 4740 -620
rect 4390 -990 4420 -810
rect 4720 -990 4740 -810
rect 4390 -1090 4740 -990
rect 2710 -1289 4740 -1090
rect 2780 -1290 4637 -1289
rect 2780 -1291 3293 -1290
rect 2780 -1349 2910 -1291
rect 2971 -1349 3099 -1291
rect 3160 -1348 3293 -1291
rect 3354 -1291 4637 -1290
rect 3354 -1348 3483 -1291
rect 3160 -1349 3483 -1348
rect 3544 -1349 3676 -1291
rect 3737 -1349 3867 -1291
rect 3928 -1349 4062 -1291
rect 4123 -1349 4252 -1291
rect 4313 -1349 4444 -1291
rect 4505 -1347 4637 -1291
rect 4698 -1347 4740 -1289
rect 4505 -1349 4740 -1347
rect 2710 -1350 4740 -1349
rect 2710 -1359 2780 -1350
rect 2910 -1359 2971 -1350
rect 3099 -1359 3160 -1350
rect 3293 -1358 3354 -1350
rect 3483 -1359 3544 -1350
rect 3676 -1359 3737 -1350
rect 3867 -1359 3928 -1350
rect 4062 -1359 4123 -1350
rect 4252 -1359 4313 -1350
rect 4444 -1359 4505 -1350
rect 4637 -1357 4698 -1350
rect 2810 -1420 2871 -1411
rect 3003 -1420 3064 -1410
rect 3194 -1420 3255 -1410
rect 3385 -1420 3446 -1412
rect 3579 -1420 3640 -1410
rect 3773 -1420 3834 -1412
rect 3962 -1420 4023 -1412
rect 4155 -1420 4216 -1412
rect 4346 -1420 4407 -1410
rect 4538 -1420 4599 -1412
rect 2690 -1421 3003 -1420
rect 2690 -1479 2810 -1421
rect 2871 -1478 3003 -1421
rect 3064 -1478 3194 -1420
rect 3255 -1422 3579 -1420
rect 3255 -1478 3385 -1422
rect 2871 -1479 3385 -1478
rect 2690 -1480 3385 -1479
rect 3446 -1478 3579 -1422
rect 3640 -1422 4346 -1420
rect 3640 -1478 3773 -1422
rect 3446 -1480 3773 -1478
rect 3834 -1480 3962 -1422
rect 4023 -1480 4155 -1422
rect 4216 -1478 4346 -1422
rect 4407 -1422 4730 -1420
rect 4407 -1478 4538 -1422
rect 4216 -1480 4538 -1478
rect 4599 -1480 4730 -1422
rect 2690 -1830 4730 -1480
rect 4330 -1950 4710 -1830
rect 4330 -2240 4360 -1950
rect 4680 -2240 4710 -1950
rect 4330 -2270 4710 -2240
use sky130_fd_pr__pfet_01v8_8DVCWJ  sky130_fd_pr__pfet_01v8_8DVCWJ_0 ~/asic/konstt-new-inv/mag
timestamp 1761646426
transform 1 0 3717 0 1 -281
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_MGS3BN  XM1
timestamp 1761646426
transform 1 0 2071 0 -1 -316
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1761646426
transform 1 0 2071 0 1 -1411
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_YTLFGX  XM4 ~/asic/konstt-new-inv/mag
timestamp 1761646426
transform 1 0 3707 0 1 -1390
box -1127 -310 1127 310
<< labels >>
flabel metal1 5200 -1000 5400 -800 0 FreeSans 256 0 0 0 out0
port 2 nsew
flabel metal1 1420 -1000 1620 -800 0 FreeSans 256 0 0 0 in0
port 3 nsew
flabel metal1 2020 -2200 2220 -2000 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 2020 200 2220 400 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
